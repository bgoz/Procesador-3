library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
entity InstructionMemory is
    Port ( rst : in  STD_LOGIC;
           address : in  STD_LOGIC_VECTOR (31 downto 0);
           imout : out  STD_LOGIC_VECTOR (31 downto 0):=(others=>'0'));
end InstructionMemory;
architecture Behavioral of InstructionMemory is
type rom_type is array (63 downto 0) of STD_LOGIC_VECTOR (31 downto 0);                 
	 signal ROM : rom_type:= (
									  "00000001000000000000000000000000",
									  "00000001000000000000000000000000",
									  "00000001000000000000000000000000",
									  "00000001000000000000000000000000",
									  "00000001000000000000000000000000",
									  "00000001000000000000000000000000",
									  "00000001000000000000000000000000",
									  "00000001000000000000000000000000",
									  "00000001000000000000000000000000",
									  "00000001000000000000000000000000",
									  "00000001000000000000000000000000",
									  "00000001000000000000000000000000",
									  "00000001000000000000000000000000",
									  "00000001000000000000000000000000",
									  "00000001000000000000000000000000",
									  "00000001000000000000000000000000",
									  "00000001000000000000000000000000",
									  "00000001000000000000000000000000",
									  "00000001000000000000000000000000",
									  "00000001000000000000000000000000",
									  "00000001000000000000000000000000",
									  "00000001000000000000000000000000",
									  "00000001000000000000000000000000",
									  "00000001000000000000000000000000",
									  "00000001000000000000000000000000",
									  "00000001000000000000000000000000",
									  "00000001000000000000000000000000",
									  "00000001000000000000000000000000",
									  "00000001000000000000000000000000",
									  "00000001000000000000000000000000",
									  "00000001000000000000000000000000",
									  "00000001000000000000000000000000",
									  "00000001000000000000000000000000",
									  "00000001000000000000000000000000",
									  "00000001000000000000000000000000",
									  "00000001000000000000000000000000",
									  "00000001000000000000000000000000",
									  "00000001000000000000000000000000",
									  "00000001000000000000000000000000",
									  "00000001000000000000000000000000",
									  "00000001000000000000000000000000",
									  "00000001000000000000000000000000",
									  "00000001000000000000000000000000",
									  "00000001000000000000000000000000",
									  "00000001000000000000000000000000",
									  "10011110000100000000000000010000", ---return o7
									  "00000001000000000000000000000000", ---nop
									  "10000001110000000010000000000011", ---jmpl 3
									  "10110010000100000010000000000100", ---mov 4 i1
									  "10110000000100000010000000000010", ---mov 2 i0 ---main
									  "00000001000000000000000000000000", ---nop
									  "10000001110000000010000000000101", ---jmpl 5
									  "10100010000101011100000000000000", ---mov %l7 %l1
									  "10101110000001000110000000000001", ---add %l7 %l1+1
									  "10100000000101011100000000000000", ---mov %l7 %l0
									  "10101110000001000000000000011000", ---add %l7 suma+%i0
									  "00000001000000000000000000000000", ---nop
									  "00000010100000000000000000001011", ---be 12 return 
									  "10000000101001000100000000011001", ---cmp %l1 %i1    ---for
									  "10100010000100000010000000000000", ---mov 0 %l1 contador
									  "10100000000100000010000000000000", ---mov 0 %l0 suma ---mult
									  "00000001000000000000000000000000", ---nop
									  "01000000000000000000000000001100", ---call 13	  
									  "00000001000000000000000000000000");
	signal rdata : std_logic_vector (31 downto 0);
begin
	rdata <= ROM(conv_integer(address));
	process (rst,address)
	begin
		  if (rst = '1') then
				imout <= ROM(conv_integer("00000000000000000000000000000000"));
		  else
				imout <= rdata;
		  end if;
	end process;
end Behavioral;							  
